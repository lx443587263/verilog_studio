//8bit 位宽加法器例化
module full_adder8(
     input [7:0]   a ,   //adder1
     input [7:0]   b ,   //adder2
      input         c ,   //input carry bit
      output        co,   //output carry bit
     output [7:0]  so   //adding result

     );

   wire [7:0]      co_temp ;
endmodule
